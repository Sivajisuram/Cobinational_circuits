`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.02.2026 17:51:24
// Design Name: 
// Module Name: half_adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module half_adder(

        input a,b,
        output  sum,carry);

   assign sum = a ^ b  ;
   assign carry = a & b; 
   
   //behavioural modelling
   /*always @ (*)begin
      
      sum = a ^ b ;
      carry = a & b ;
      end */
endmodule
